module carry_lookahead(input [15:0] A,B, input cin, output logic [15:0] sum, output logic cout);
